`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:51:07 05/28/2016 
// Design Name: 
// Module Name:    pic_ram 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pic_ram(
	clk,
	rst,
	addr,
	data_out
    );
	input clk;
	input rst;
	input [9:0] addr;
	output reg [7:0] data_out;
	
	reg [7:0] pic [0:783];
	reg cnt;
	
	always @ (posedge clk) begin
		if (rst) begin
			//picture
		  //addr <= 10'd0;
		  data_out <= pic[0];
        pic[ 0 ] <= 8'd 0 ;
        pic[ 1 ] <= 8'd 0 ;
        pic[ 2 ] <= 8'd 0 ;
        pic[ 3 ] <= 8'd 0 ;
        pic[ 4 ] <= 8'd 0 ;
        pic[ 5 ] <= 8'd 0 ;
        pic[ 6 ] <= 8'd 0 ;
        pic[ 7 ] <= 8'd 0 ;
        pic[ 8 ] <= 8'd 0 ;
        pic[ 9 ] <= 8'd 0 ;
        pic[ 10 ] <= 8'd 0 ;
        pic[ 11 ] <= 8'd 0 ;
        pic[ 12 ] <= 8'd 0 ;
        pic[ 13 ] <= 8'd 0 ;
        pic[ 14 ] <= 8'd 0 ;
        pic[ 15 ] <= 8'd 0 ;
        pic[ 16 ] <= 8'd 0 ;
        pic[ 17 ] <= 8'd 0 ;
        pic[ 18 ] <= 8'd 0 ;
        pic[ 19 ] <= 8'd 0 ;
        pic[ 20 ] <= 8'd 0 ;
        pic[ 21 ] <= 8'd 0 ;
        pic[ 22 ] <= 8'd 0 ;
        pic[ 23 ] <= 8'd 0 ;
        pic[ 24 ] <= 8'd 0 ;
        pic[ 25 ] <= 8'd 0 ;
        pic[ 26 ] <= 8'd 0 ;
        pic[ 27 ] <= 8'd 0 ;
        pic[ 28 ] <= 8'd 0 ;
        pic[ 29 ] <= 8'd 0 ;
        pic[ 30 ] <= 8'd 0 ;
        pic[ 31 ] <= 8'd 0 ;
        pic[ 32 ] <= 8'd 0 ;
        pic[ 33 ] <= 8'd 0 ;
        pic[ 34 ] <= 8'd 0 ;
        pic[ 35 ] <= 8'd 0 ;
        pic[ 36 ] <= 8'd 0 ;
        pic[ 37 ] <= 8'd 0 ;
        pic[ 38 ] <= 8'd 0 ;
        pic[ 39 ] <= 8'd 0 ;
        pic[ 40 ] <= 8'd 0 ;
        pic[ 41 ] <= 8'd 0 ;
        pic[ 42 ] <= 8'd 0 ;
        pic[ 43 ] <= 8'd 0 ;
        pic[ 44 ] <= 8'd 0 ;
        pic[ 45 ] <= 8'd 0 ;
        pic[ 46 ] <= 8'd 0 ;
        pic[ 47 ] <= 8'd 0 ;
        pic[ 48 ] <= 8'd 0 ;
        pic[ 49 ] <= 8'd 0 ;
        pic[ 50 ] <= 8'd 0 ;
        pic[ 51 ] <= 8'd 0 ;
        pic[ 52 ] <= 8'd 0 ;
        pic[ 53 ] <= 8'd 0 ;
        pic[ 54 ] <= 8'd 0 ;
        pic[ 55 ] <= 8'd 0 ;
        pic[ 56 ] <= 8'd 0 ;
        pic[ 57 ] <= 8'd 0 ;
        pic[ 58 ] <= 8'd 0 ;
        pic[ 59 ] <= 8'd 0 ;
        pic[ 60 ] <= 8'd 0 ;
        pic[ 61 ] <= 8'd 0 ;
        pic[ 62 ] <= 8'd 0 ;
        pic[ 63 ] <= 8'd 0 ;
        pic[ 64 ] <= 8'd 0 ;
        pic[ 65 ] <= 8'd 0 ;
        pic[ 66 ] <= 8'd 0 ;
        pic[ 67 ] <= 8'd 0 ;
        pic[ 68 ] <= 8'd 0 ;
        pic[ 69 ] <= 8'd 0 ;
        pic[ 70 ] <= 8'd 0 ;
        pic[ 71 ] <= 8'd 0 ;
        pic[ 72 ] <= 8'd 0 ;
        pic[ 73 ] <= 8'd 0 ;
        pic[ 74 ] <= 8'd 0 ;
        pic[ 75 ] <= 8'd 0 ;
        pic[ 76 ] <= 8'd 0 ;
        pic[ 77 ] <= 8'd 0 ;
        pic[ 78 ] <= 8'd 0 ;
        pic[ 79 ] <= 8'd 0 ;
        pic[ 80 ] <= 8'd 0 ;
        pic[ 81 ] <= 8'd 0 ;
        pic[ 82 ] <= 8'd 0 ;
        pic[ 83 ] <= 8'd 0 ;
        pic[ 84 ] <= 8'd 0 ;
        pic[ 85 ] <= 8'd 0 ;
        pic[ 86 ] <= 8'd 0 ;
        pic[ 87 ] <= 8'd 0 ;
        pic[ 88 ] <= 8'd 0 ;
        pic[ 89 ] <= 8'd 0 ;
        pic[ 90 ] <= 8'd 0 ;
        pic[ 91 ] <= 8'd 0 ;
        pic[ 92 ] <= 8'd 0 ;
        pic[ 93 ] <= 8'd 0 ;
        pic[ 94 ] <= 8'd 0 ;
        pic[ 95 ] <= 8'd 0 ;
        pic[ 96 ] <= 8'd 0 ;
        pic[ 97 ] <= 8'd 0 ;
        pic[ 98 ] <= 8'd 0 ;
        pic[ 99 ] <= 8'd 0 ;
        pic[ 100 ] <= 8'd 0 ;
        pic[ 101 ] <= 8'd 0 ;
        pic[ 102 ] <= 8'd 0 ;
        pic[ 103 ] <= 8'd 0 ;
        pic[ 104 ] <= 8'd 0 ;
        pic[ 105 ] <= 8'd 0 ;
        pic[ 106 ] <= 8'd 0 ;
        pic[ 107 ] <= 8'd 0 ;
        pic[ 108 ] <= 8'd 0 ;
        pic[ 109 ] <= 8'd 0 ;
        pic[ 110 ] <= 8'd 0 ;
        pic[ 111 ] <= 8'd 0 ;
        pic[ 112 ] <= 8'd 0 ;
        pic[ 113 ] <= 8'd 0 ;
        pic[ 114 ] <= 8'd 0 ;
        pic[ 115 ] <= 8'd 0 ;
        pic[ 116 ] <= 8'd 0 ;
        pic[ 117 ] <= 8'd 0 ;
        pic[ 118 ] <= 8'd 0 ;
        pic[ 119 ] <= 8'd 0 ;
        pic[ 120 ] <= 8'd 0 ;
        pic[ 121 ] <= 8'd 0 ;
        pic[ 122 ] <= 8'd 0 ;
        pic[ 123 ] <= 8'd 0 ;
        pic[ 124 ] <= 8'd 0 ;
        pic[ 125 ] <= 8'd 0 ;
        pic[ 126 ] <= 8'd 0 ;
        pic[ 127 ] <= 8'd 0 ;
        pic[ 128 ] <= 8'd 38 ;
        pic[ 129 ] <= 8'd 254 ;
        pic[ 130 ] <= 8'd 109 ;
        pic[ 131 ] <= 8'd 0 ;
        pic[ 132 ] <= 8'd 0 ;
        pic[ 133 ] <= 8'd 0 ;
        pic[ 134 ] <= 8'd 0 ;
        pic[ 135 ] <= 8'd 0 ;
        pic[ 136 ] <= 8'd 0 ;
        pic[ 137 ] <= 8'd 0 ;
        pic[ 138 ] <= 8'd 0 ;
        pic[ 139 ] <= 8'd 0 ;
        pic[ 140 ] <= 8'd 0 ;
        pic[ 141 ] <= 8'd 0 ;
        pic[ 142 ] <= 8'd 0 ;
        pic[ 143 ] <= 8'd 0 ;
        pic[ 144 ] <= 8'd 0 ;
        pic[ 145 ] <= 8'd 0 ;
        pic[ 146 ] <= 8'd 0 ;
        pic[ 147 ] <= 8'd 0 ;
        pic[ 148 ] <= 8'd 0 ;
        pic[ 149 ] <= 8'd 0 ;
        pic[ 150 ] <= 8'd 0 ;
        pic[ 151 ] <= 8'd 0 ;
        pic[ 152 ] <= 8'd 0 ;
        pic[ 153 ] <= 8'd 0 ;
        pic[ 154 ] <= 8'd 0 ;
        pic[ 155 ] <= 8'd 0 ;
        pic[ 156 ] <= 8'd 87 ;
        pic[ 157 ] <= 8'd 252 ;
        pic[ 158 ] <= 8'd 82 ;
        pic[ 159 ] <= 8'd 0 ;
        pic[ 160 ] <= 8'd 0 ;
        pic[ 161 ] <= 8'd 0 ;
        pic[ 162 ] <= 8'd 0 ;
        pic[ 163 ] <= 8'd 0 ;
        pic[ 164 ] <= 8'd 0 ;
        pic[ 165 ] <= 8'd 0 ;
        pic[ 166 ] <= 8'd 0 ;
        pic[ 167 ] <= 8'd 0 ;
        pic[ 168 ] <= 8'd 0 ;
        pic[ 169 ] <= 8'd 0 ;
        pic[ 170 ] <= 8'd 0 ;
        pic[ 171 ] <= 8'd 0 ;
        pic[ 172 ] <= 8'd 0 ;
        pic[ 173 ] <= 8'd 0 ;
        pic[ 174 ] <= 8'd 0 ;
        pic[ 175 ] <= 8'd 0 ;
        pic[ 176 ] <= 8'd 0 ;
        pic[ 177 ] <= 8'd 0 ;
        pic[ 178 ] <= 8'd 0 ;
        pic[ 179 ] <= 8'd 0 ;
        pic[ 180 ] <= 8'd 0 ;
        pic[ 181 ] <= 8'd 0 ;
        pic[ 182 ] <= 8'd 0 ;
        pic[ 183 ] <= 8'd 0 ;
        pic[ 184 ] <= 8'd 135 ;
        pic[ 185 ] <= 8'd 241 ;
        pic[ 186 ] <= 8'd 0 ;
        pic[ 187 ] <= 8'd 0 ;
        pic[ 188 ] <= 8'd 0 ;
        pic[ 189 ] <= 8'd 0 ;
        pic[ 190 ] <= 8'd 0 ;
        pic[ 191 ] <= 8'd 0 ;
        pic[ 192 ] <= 8'd 0 ;
        pic[ 193 ] <= 8'd 0 ;
        pic[ 194 ] <= 8'd 0 ;
        pic[ 195 ] <= 8'd 0 ;
        pic[ 196 ] <= 8'd 0 ;
        pic[ 197 ] <= 8'd 0 ;
        pic[ 198 ] <= 8'd 0 ;
        pic[ 199 ] <= 8'd 0 ;
        pic[ 200 ] <= 8'd 0 ;
        pic[ 201 ] <= 8'd 0 ;
        pic[ 202 ] <= 8'd 0 ;
        pic[ 203 ] <= 8'd 0 ;
        pic[ 204 ] <= 8'd 0 ;
        pic[ 205 ] <= 8'd 0 ;
        pic[ 206 ] <= 8'd 0 ;
        pic[ 207 ] <= 8'd 0 ;
        pic[ 208 ] <= 8'd 0 ;
        pic[ 209 ] <= 8'd 0 ;
        pic[ 210 ] <= 8'd 0 ;
        pic[ 211 ] <= 8'd 45 ;
        pic[ 212 ] <= 8'd 244 ;
        pic[ 213 ] <= 8'd 150 ;
        pic[ 214 ] <= 8'd 0 ;
        pic[ 215 ] <= 8'd 0 ;
        pic[ 216 ] <= 8'd 0 ;
        pic[ 217 ] <= 8'd 0 ;
        pic[ 218 ] <= 8'd 0 ;
        pic[ 219 ] <= 8'd 0 ;
        pic[ 220 ] <= 8'd 0 ;
        pic[ 221 ] <= 8'd 0 ;
        pic[ 222 ] <= 8'd 0 ;
        pic[ 223 ] <= 8'd 0 ;
        pic[ 224 ] <= 8'd 0 ;
        pic[ 225 ] <= 8'd 0 ;
        pic[ 226 ] <= 8'd 0 ;
        pic[ 227 ] <= 8'd 0 ;
        pic[ 228 ] <= 8'd 0 ;
        pic[ 229 ] <= 8'd 0 ;
        pic[ 230 ] <= 8'd 0 ;
        pic[ 231 ] <= 8'd 0 ;
        pic[ 232 ] <= 8'd 0 ;
        pic[ 233 ] <= 8'd 0 ;
        pic[ 234 ] <= 8'd 0 ;
        pic[ 235 ] <= 8'd 0 ;
        pic[ 236 ] <= 8'd 0 ;
        pic[ 237 ] <= 8'd 0 ;
        pic[ 238 ] <= 8'd 0 ;
        pic[ 239 ] <= 8'd 84 ;
        pic[ 240 ] <= 8'd 254 ;
        pic[ 241 ] <= 8'd 63 ;
        pic[ 242 ] <= 8'd 0 ;
        pic[ 243 ] <= 8'd 0 ;
        pic[ 244 ] <= 8'd 0 ;
        pic[ 245 ] <= 8'd 0 ;
        pic[ 246 ] <= 8'd 0 ;
        pic[ 247 ] <= 8'd 0 ;
        pic[ 248 ] <= 8'd 0 ;
        pic[ 249 ] <= 8'd 0 ;
        pic[ 250 ] <= 8'd 0 ;
        pic[ 251 ] <= 8'd 0 ;
        pic[ 252 ] <= 8'd 0 ;
        pic[ 253 ] <= 8'd 0 ;
        pic[ 254 ] <= 8'd 0 ;
        pic[ 255 ] <= 8'd 0 ;
        pic[ 256 ] <= 8'd 0 ;
        pic[ 257 ] <= 8'd 0 ;
        pic[ 258 ] <= 8'd 0 ;
        pic[ 259 ] <= 8'd 0 ;
        pic[ 260 ] <= 8'd 0 ;
        pic[ 261 ] <= 8'd 0 ;
        pic[ 262 ] <= 8'd 0 ;
        pic[ 263 ] <= 8'd 0 ;
        pic[ 264 ] <= 8'd 0 ;
        pic[ 265 ] <= 8'd 0 ;
        pic[ 266 ] <= 8'd 0 ;
        pic[ 267 ] <= 8'd 202 ;
        pic[ 268 ] <= 8'd 223 ;
        pic[ 269 ] <= 8'd 11 ;
        pic[ 270 ] <= 8'd 0 ;
        pic[ 271 ] <= 8'd 0 ;
        pic[ 272 ] <= 8'd 0 ;
        pic[ 273 ] <= 8'd 0 ;
        pic[ 274 ] <= 8'd 0 ;
        pic[ 275 ] <= 8'd 0 ;
        pic[ 276 ] <= 8'd 0 ;
        pic[ 277 ] <= 8'd 0 ;
        pic[ 278 ] <= 8'd 0 ;
        pic[ 279 ] <= 8'd 0 ;
        pic[ 280 ] <= 8'd 0 ;
        pic[ 281 ] <= 8'd 0 ;
        pic[ 282 ] <= 8'd 0 ;
        pic[ 283 ] <= 8'd 0 ;
        pic[ 284 ] <= 8'd 0 ;
        pic[ 285 ] <= 8'd 0 ;
        pic[ 286 ] <= 8'd 0 ;
        pic[ 287 ] <= 8'd 0 ;
        pic[ 288 ] <= 8'd 0 ;
        pic[ 289 ] <= 8'd 0 ;
        pic[ 290 ] <= 8'd 0 ;
        pic[ 291 ] <= 8'd 0 ;
        pic[ 292 ] <= 8'd 0 ;
        pic[ 293 ] <= 8'd 0 ;
        pic[ 294 ] <= 8'd 32 ;
        pic[ 295 ] <= 8'd 254 ;
        pic[ 296 ] <= 8'd 216 ;
        pic[ 297 ] <= 8'd 0 ;
        pic[ 298 ] <= 8'd 0 ;
        pic[ 299 ] <= 8'd 0 ;
        pic[ 300 ] <= 8'd 0 ;
        pic[ 301 ] <= 8'd 0 ;
        pic[ 302 ] <= 8'd 0 ;
        pic[ 303 ] <= 8'd 0 ;
        pic[ 304 ] <= 8'd 0 ;
        pic[ 305 ] <= 8'd 0 ;
        pic[ 306 ] <= 8'd 0 ;
        pic[ 307 ] <= 8'd 0 ;
        pic[ 308 ] <= 8'd 0 ;
        pic[ 309 ] <= 8'd 0 ;
        pic[ 310 ] <= 8'd 0 ;
        pic[ 311 ] <= 8'd 0 ;
        pic[ 312 ] <= 8'd 0 ;
        pic[ 313 ] <= 8'd 0 ;
        pic[ 314 ] <= 8'd 0 ;
        pic[ 315 ] <= 8'd 0 ;
        pic[ 316 ] <= 8'd 0 ;
        pic[ 317 ] <= 8'd 0 ;
        pic[ 318 ] <= 8'd 0 ;
        pic[ 319 ] <= 8'd 0 ;
        pic[ 320 ] <= 8'd 0 ;
        pic[ 321 ] <= 8'd 0 ;
        pic[ 322 ] <= 8'd 95 ;
        pic[ 323 ] <= 8'd 254 ;
        pic[ 324 ] <= 8'd 195 ;
        pic[ 325 ] <= 8'd 0 ;
        pic[ 326 ] <= 8'd 0 ;
        pic[ 327 ] <= 8'd 0 ;
        pic[ 328 ] <= 8'd 0 ;
        pic[ 329 ] <= 8'd 0 ;
        pic[ 330 ] <= 8'd 0 ;
        pic[ 331 ] <= 8'd 0 ;
        pic[ 332 ] <= 8'd 0 ;
        pic[ 333 ] <= 8'd 0 ;
        pic[ 334 ] <= 8'd 0 ;
        pic[ 335 ] <= 8'd 0 ;
        pic[ 336 ] <= 8'd 0 ;
        pic[ 337 ] <= 8'd 0 ;
        pic[ 338 ] <= 8'd 0 ;
        pic[ 339 ] <= 8'd 0 ;
        pic[ 340 ] <= 8'd 0 ;
        pic[ 341 ] <= 8'd 0 ;
        pic[ 342 ] <= 8'd 0 ;
        pic[ 343 ] <= 8'd 0 ;
        pic[ 344 ] <= 8'd 0 ;
        pic[ 345 ] <= 8'd 0 ;
        pic[ 346 ] <= 8'd 0 ;
        pic[ 347 ] <= 8'd 0 ;
        pic[ 348 ] <= 8'd 0 ;
        pic[ 349 ] <= 8'd 0 ;
        pic[ 350 ] <= 8'd 140 ;
        pic[ 351 ] <= 8'd 254 ;
        pic[ 352 ] <= 8'd 77 ;
        pic[ 353 ] <= 8'd 0 ;
        pic[ 354 ] <= 8'd 0 ;
        pic[ 355 ] <= 8'd 0 ;
        pic[ 356 ] <= 8'd 0 ;
        pic[ 357 ] <= 8'd 0 ;
        pic[ 358 ] <= 8'd 0 ;
        pic[ 359 ] <= 8'd 0 ;
        pic[ 360 ] <= 8'd 0 ;
        pic[ 361 ] <= 8'd 0 ;
        pic[ 362 ] <= 8'd 0 ;
        pic[ 363 ] <= 8'd 0 ;
        pic[ 364 ] <= 8'd 0 ;
        pic[ 365 ] <= 8'd 0 ;
        pic[ 366 ] <= 8'd 0 ;
        pic[ 367 ] <= 8'd 0 ;
        pic[ 368 ] <= 8'd 0 ;
        pic[ 369 ] <= 8'd 0 ;
        pic[ 370 ] <= 8'd 0 ;
        pic[ 371 ] <= 8'd 0 ;
        pic[ 372 ] <= 8'd 0 ;
        pic[ 373 ] <= 8'd 0 ;
        pic[ 374 ] <= 8'd 0 ;
        pic[ 375 ] <= 8'd 0 ;
        pic[ 376 ] <= 8'd 0 ;
        pic[ 377 ] <= 8'd 57 ;
        pic[ 378 ] <= 8'd 237 ;
        pic[ 379 ] <= 8'd 205 ;
        pic[ 380 ] <= 8'd 8 ;
        pic[ 381 ] <= 8'd 0 ;
        pic[ 382 ] <= 8'd 0 ;
        pic[ 383 ] <= 8'd 0 ;
        pic[ 384 ] <= 8'd 0 ;
        pic[ 385 ] <= 8'd 0 ;
        pic[ 386 ] <= 8'd 0 ;
        pic[ 387 ] <= 8'd 0 ;
        pic[ 388 ] <= 8'd 0 ;
        pic[ 389 ] <= 8'd 0 ;
        pic[ 390 ] <= 8'd 0 ;
        pic[ 391 ] <= 8'd 0 ;
        pic[ 392 ] <= 8'd 0 ;
        pic[ 393 ] <= 8'd 0 ;
        pic[ 394 ] <= 8'd 0 ;
        pic[ 395 ] <= 8'd 0 ;
        pic[ 396 ] <= 8'd 0 ;
        pic[ 397 ] <= 8'd 0 ;
        pic[ 398 ] <= 8'd 0 ;
        pic[ 399 ] <= 8'd 0 ;
        pic[ 400 ] <= 8'd 0 ;
        pic[ 401 ] <= 8'd 0 ;
        pic[ 402 ] <= 8'd 0 ;
        pic[ 403 ] <= 8'd 0 ;
        pic[ 404 ] <= 8'd 0 ;
        pic[ 405 ] <= 8'd 124 ;
        pic[ 406 ] <= 8'd 255 ;
        pic[ 407 ] <= 8'd 165 ;
        pic[ 408 ] <= 8'd 0 ;
        pic[ 409 ] <= 8'd 0 ;
        pic[ 410 ] <= 8'd 0 ;
        pic[ 411 ] <= 8'd 0 ;
        pic[ 412 ] <= 8'd 0 ;
        pic[ 413 ] <= 8'd 0 ;
        pic[ 414 ] <= 8'd 0 ;
        pic[ 415 ] <= 8'd 0 ;
        pic[ 416 ] <= 8'd 0 ;
        pic[ 417 ] <= 8'd 0 ;
        pic[ 418 ] <= 8'd 0 ;
        pic[ 419 ] <= 8'd 0 ;
        pic[ 420 ] <= 8'd 0 ;
        pic[ 421 ] <= 8'd 0 ;
        pic[ 422 ] <= 8'd 0 ;
        pic[ 423 ] <= 8'd 0 ;
        pic[ 424 ] <= 8'd 0 ;
        pic[ 425 ] <= 8'd 0 ;
        pic[ 426 ] <= 8'd 0 ;
        pic[ 427 ] <= 8'd 0 ;
        pic[ 428 ] <= 8'd 0 ;
        pic[ 429 ] <= 8'd 0 ;
        pic[ 430 ] <= 8'd 0 ;
        pic[ 431 ] <= 8'd 0 ;
        pic[ 432 ] <= 8'd 0 ;
        pic[ 433 ] <= 8'd 171 ;
        pic[ 434 ] <= 8'd 254 ;
        pic[ 435 ] <= 8'd 81 ;
        pic[ 436 ] <= 8'd 0 ;
        pic[ 437 ] <= 8'd 0 ;
        pic[ 438 ] <= 8'd 0 ;
        pic[ 439 ] <= 8'd 0 ;
        pic[ 440 ] <= 8'd 0 ;
        pic[ 441 ] <= 8'd 0 ;
        pic[ 442 ] <= 8'd 0 ;
        pic[ 443 ] <= 8'd 0 ;
        pic[ 444 ] <= 8'd 0 ;
        pic[ 445 ] <= 8'd 0 ;
        pic[ 446 ] <= 8'd 0 ;
        pic[ 447 ] <= 8'd 0 ;
        pic[ 448 ] <= 8'd 0 ;
        pic[ 449 ] <= 8'd 0 ;
        pic[ 450 ] <= 8'd 0 ;
        pic[ 451 ] <= 8'd 0 ;
        pic[ 452 ] <= 8'd 0 ;
        pic[ 453 ] <= 8'd 0 ;
        pic[ 454 ] <= 8'd 0 ;
        pic[ 455 ] <= 8'd 0 ;
        pic[ 456 ] <= 8'd 0 ;
        pic[ 457 ] <= 8'd 0 ;
        pic[ 458 ] <= 8'd 0 ;
        pic[ 459 ] <= 8'd 0 ;
        pic[ 460 ] <= 8'd 24 ;
        pic[ 461 ] <= 8'd 232 ;
        pic[ 462 ] <= 8'd 215 ;
        pic[ 463 ] <= 8'd 0 ;
        pic[ 464 ] <= 8'd 0 ;
        pic[ 465 ] <= 8'd 0 ;
        pic[ 466 ] <= 8'd 0 ;
        pic[ 467 ] <= 8'd 0 ;
        pic[ 468 ] <= 8'd 0 ;
        pic[ 469 ] <= 8'd 0 ;
        pic[ 470 ] <= 8'd 0 ;
        pic[ 471 ] <= 8'd 0 ;
        pic[ 472 ] <= 8'd 0 ;
        pic[ 473 ] <= 8'd 0 ;
        pic[ 474 ] <= 8'd 0 ;
        pic[ 475 ] <= 8'd 0 ;
        pic[ 476 ] <= 8'd 0 ;
        pic[ 477 ] <= 8'd 0 ;
        pic[ 478 ] <= 8'd 0 ;
        pic[ 479 ] <= 8'd 0 ;
        pic[ 480 ] <= 8'd 0 ;
        pic[ 481 ] <= 8'd 0 ;
        pic[ 482 ] <= 8'd 0 ;
        pic[ 483 ] <= 8'd 0 ;
        pic[ 484 ] <= 8'd 0 ;
        pic[ 485 ] <= 8'd 0 ;
        pic[ 486 ] <= 8'd 0 ;
        pic[ 487 ] <= 8'd 0 ;
        pic[ 488 ] <= 8'd 120 ;
        pic[ 489 ] <= 8'd 254 ;
        pic[ 490 ] <= 8'd 159 ;
        pic[ 491 ] <= 8'd 0 ;
        pic[ 492 ] <= 8'd 0 ;
        pic[ 493 ] <= 8'd 0 ;
        pic[ 494 ] <= 8'd 0 ;
        pic[ 495 ] <= 8'd 0 ;
        pic[ 496 ] <= 8'd 0 ;
        pic[ 497 ] <= 8'd 0 ;
        pic[ 498 ] <= 8'd 0 ;
        pic[ 499 ] <= 8'd 0 ;
        pic[ 500 ] <= 8'd 0 ;
        pic[ 501 ] <= 8'd 0 ;
        pic[ 502 ] <= 8'd 0 ;
        pic[ 503 ] <= 8'd 0 ;
        pic[ 504 ] <= 8'd 0 ;
        pic[ 505 ] <= 8'd 0 ;
        pic[ 506 ] <= 8'd 0 ;
        pic[ 507 ] <= 8'd 0 ;
        pic[ 508 ] <= 8'd 0 ;
        pic[ 509 ] <= 8'd 0 ;
        pic[ 510 ] <= 8'd 0 ;
        pic[ 511 ] <= 8'd 0 ;
        pic[ 512 ] <= 8'd 0 ;
        pic[ 513 ] <= 8'd 0 ;
        pic[ 514 ] <= 8'd 0 ;
        pic[ 515 ] <= 8'd 0 ;
        pic[ 516 ] <= 8'd 151 ;
        pic[ 517 ] <= 8'd 254 ;
        pic[ 518 ] <= 8'd 142 ;
        pic[ 519 ] <= 8'd 0 ;
        pic[ 520 ] <= 8'd 0 ;
        pic[ 521 ] <= 8'd 0 ;
        pic[ 522 ] <= 8'd 0 ;
        pic[ 523 ] <= 8'd 0 ;
        pic[ 524 ] <= 8'd 0 ;
        pic[ 525 ] <= 8'd 0 ;
        pic[ 526 ] <= 8'd 0 ;
        pic[ 527 ] <= 8'd 0 ;
        pic[ 528 ] <= 8'd 0 ;
        pic[ 529 ] <= 8'd 0 ;
        pic[ 530 ] <= 8'd 0 ;
        pic[ 531 ] <= 8'd 0 ;
        pic[ 532 ] <= 8'd 0 ;
        pic[ 533 ] <= 8'd 0 ;
        pic[ 534 ] <= 8'd 0 ;
        pic[ 535 ] <= 8'd 0 ;
        pic[ 536 ] <= 8'd 0 ;
        pic[ 537 ] <= 8'd 0 ;
        pic[ 538 ] <= 8'd 0 ;
        pic[ 539 ] <= 8'd 0 ;
        pic[ 540 ] <= 8'd 0 ;
        pic[ 541 ] <= 8'd 0 ;
        pic[ 542 ] <= 8'd 0 ;
        pic[ 543 ] <= 8'd 0 ;
        pic[ 544 ] <= 8'd 228 ;
        pic[ 545 ] <= 8'd 254 ;
        pic[ 546 ] <= 8'd 66 ;
        pic[ 547 ] <= 8'd 0 ;
        pic[ 548 ] <= 8'd 0 ;
        pic[ 549 ] <= 8'd 0 ;
        pic[ 550 ] <= 8'd 0 ;
        pic[ 551 ] <= 8'd 0 ;
        pic[ 552 ] <= 8'd 0 ;
        pic[ 553 ] <= 8'd 0 ;
        pic[ 554 ] <= 8'd 0 ;
        pic[ 555 ] <= 8'd 0 ;
        pic[ 556 ] <= 8'd 0 ;
        pic[ 557 ] <= 8'd 0 ;
        pic[ 558 ] <= 8'd 0 ;
        pic[ 559 ] <= 8'd 0 ;
        pic[ 560 ] <= 8'd 0 ;
        pic[ 561 ] <= 8'd 0 ;
        pic[ 562 ] <= 8'd 0 ;
        pic[ 563 ] <= 8'd 0 ;
        pic[ 564 ] <= 8'd 0 ;
        pic[ 565 ] <= 8'd 0 ;
        pic[ 566 ] <= 8'd 0 ;
        pic[ 567 ] <= 8'd 0 ;
        pic[ 568 ] <= 8'd 0 ;
        pic[ 569 ] <= 8'd 0 ;
        pic[ 570 ] <= 8'd 0 ;
        pic[ 571 ] <= 8'd 61 ;
        pic[ 572 ] <= 8'd 251 ;
        pic[ 573 ] <= 8'd 254 ;
        pic[ 574 ] <= 8'd 66 ;
        pic[ 575 ] <= 8'd 0 ;
        pic[ 576 ] <= 8'd 0 ;
        pic[ 577 ] <= 8'd 0 ;
        pic[ 578 ] <= 8'd 0 ;
        pic[ 579 ] <= 8'd 0 ;
        pic[ 580 ] <= 8'd 0 ;
        pic[ 581 ] <= 8'd 0 ;
        pic[ 582 ] <= 8'd 0 ;
        pic[ 583 ] <= 8'd 0 ;
        pic[ 584 ] <= 8'd 0 ;
        pic[ 585 ] <= 8'd 0 ;
        pic[ 586 ] <= 8'd 0 ;
        pic[ 587 ] <= 8'd 0 ;
        pic[ 588 ] <= 8'd 0 ;
        pic[ 589 ] <= 8'd 0 ;
        pic[ 590 ] <= 8'd 0 ;
        pic[ 591 ] <= 8'd 0 ;
        pic[ 592 ] <= 8'd 0 ;
        pic[ 593 ] <= 8'd 0 ;
        pic[ 594 ] <= 8'd 0 ;
        pic[ 595 ] <= 8'd 0 ;
        pic[ 596 ] <= 8'd 0 ;
        pic[ 597 ] <= 8'd 0 ;
        pic[ 598 ] <= 8'd 0 ;
        pic[ 599 ] <= 8'd 141 ;
        pic[ 600 ] <= 8'd 254 ;
        pic[ 601 ] <= 8'd 205 ;
        pic[ 602 ] <= 8'd 3 ;
        pic[ 603 ] <= 8'd 0 ;
        pic[ 604 ] <= 8'd 0 ;
        pic[ 605 ] <= 8'd 0 ;
        pic[ 606 ] <= 8'd 0 ;
        pic[ 607 ] <= 8'd 0 ;
        pic[ 608 ] <= 8'd 0 ;
        pic[ 609 ] <= 8'd 0 ;
        pic[ 610 ] <= 8'd 0 ;
        pic[ 611 ] <= 8'd 0 ;
        pic[ 612 ] <= 8'd 0 ;
        pic[ 613 ] <= 8'd 0 ;
        pic[ 614 ] <= 8'd 0 ;
        pic[ 615 ] <= 8'd 0 ;
        pic[ 616 ] <= 8'd 0 ;
        pic[ 617 ] <= 8'd 0 ;
        pic[ 618 ] <= 8'd 0 ;
        pic[ 619 ] <= 8'd 0 ;
        pic[ 620 ] <= 8'd 0 ;
        pic[ 621 ] <= 8'd 0 ;
        pic[ 622 ] <= 8'd 0 ;
        pic[ 623 ] <= 8'd 0 ;
        pic[ 624 ] <= 8'd 0 ;
        pic[ 625 ] <= 8'd 0 ;
        pic[ 626 ] <= 8'd 10 ;
        pic[ 627 ] <= 8'd 215 ;
        pic[ 628 ] <= 8'd 254 ;
        pic[ 629 ] <= 8'd 121 ;
        pic[ 630 ] <= 8'd 0 ;
        pic[ 631 ] <= 8'd 0 ;
        pic[ 632 ] <= 8'd 0 ;
        pic[ 633 ] <= 8'd 0 ;
        pic[ 634 ] <= 8'd 0 ;
        pic[ 635 ] <= 8'd 0 ;
        pic[ 636 ] <= 8'd 0 ;
        pic[ 637 ] <= 8'd 0 ;
        pic[ 638 ] <= 8'd 0 ;
        pic[ 639 ] <= 8'd 0 ;
        pic[ 640 ] <= 8'd 0 ;
        pic[ 641 ] <= 8'd 0 ;
        pic[ 642 ] <= 8'd 0 ;
        pic[ 643 ] <= 8'd 0 ;
        pic[ 644 ] <= 8'd 0 ;
        pic[ 645 ] <= 8'd 0 ;
        pic[ 646 ] <= 8'd 0 ;
        pic[ 647 ] <= 8'd 0 ;
        pic[ 648 ] <= 8'd 0 ;
        pic[ 649 ] <= 8'd 0 ;
        pic[ 650 ] <= 8'd 0 ;
        pic[ 651 ] <= 8'd 0 ;
        pic[ 652 ] <= 8'd 0 ;
        pic[ 653 ] <= 8'd 0 ;
        pic[ 654 ] <= 8'd 5 ;
        pic[ 655 ] <= 8'd 198 ;
        pic[ 656 ] <= 8'd 176 ;
        pic[ 657 ] <= 8'd 10 ;
        pic[ 658 ] <= 8'd 0 ;
        pic[ 659 ] <= 8'd 0 ;
        pic[ 660 ] <= 8'd 0 ;
        pic[ 661 ] <= 8'd 0 ;
        pic[ 662 ] <= 8'd 0 ;
        pic[ 663 ] <= 8'd 0 ;
        pic[ 664 ] <= 8'd 0 ;
        pic[ 665 ] <= 8'd 0 ;
        pic[ 666 ] <= 8'd 0 ;
        pic[ 667 ] <= 8'd 0 ;
        pic[ 668 ] <= 8'd 0 ;
        pic[ 669 ] <= 8'd 0 ;
        pic[ 670 ] <= 8'd 0 ;
        pic[ 671 ] <= 8'd 0 ;
        pic[ 672 ] <= 8'd 0 ;
        pic[ 673 ] <= 8'd 0 ;
        pic[ 674 ] <= 8'd 0 ;
        pic[ 675 ] <= 8'd 0 ;
        pic[ 676 ] <= 8'd 0 ;
        pic[ 677 ] <= 8'd 0 ;
        pic[ 678 ] <= 8'd 0 ;
        pic[ 679 ] <= 8'd 0 ;
        pic[ 680 ] <= 8'd 0 ;
        pic[ 681 ] <= 8'd 0 ;
        pic[ 682 ] <= 8'd 0 ;
        pic[ 683 ] <= 8'd 0 ;
        pic[ 684 ] <= 8'd 0 ;
        pic[ 685 ] <= 8'd 0 ;
        pic[ 686 ] <= 8'd 0 ;
        pic[ 687 ] <= 8'd 0 ;
        pic[ 688 ] <= 8'd 0 ;
        pic[ 689 ] <= 8'd 0 ;
        pic[ 690 ] <= 8'd 0 ;
        pic[ 691 ] <= 8'd 0 ;
        pic[ 692 ] <= 8'd 0 ;
        pic[ 693 ] <= 8'd 0 ;
        pic[ 694 ] <= 8'd 0 ;
        pic[ 695 ] <= 8'd 0 ;
        pic[ 696 ] <= 8'd 0 ;
        pic[ 697 ] <= 8'd 0 ;
        pic[ 698 ] <= 8'd 0 ;
        pic[ 699 ] <= 8'd 0 ;
        pic[ 700 ] <= 8'd 0 ;
        pic[ 701 ] <= 8'd 0 ;
        pic[ 702 ] <= 8'd 0 ;
        pic[ 703 ] <= 8'd 0 ;
        pic[ 704 ] <= 8'd 0 ;
        pic[ 705 ] <= 8'd 0 ;
        pic[ 706 ] <= 8'd 0 ;
        pic[ 707 ] <= 8'd 0 ;
        pic[ 708 ] <= 8'd 0 ;
        pic[ 709 ] <= 8'd 0 ;
        pic[ 710 ] <= 8'd 0 ;
        pic[ 711 ] <= 8'd 0 ;
        pic[ 712 ] <= 8'd 0 ;
        pic[ 713 ] <= 8'd 0 ;
        pic[ 714 ] <= 8'd 0 ;
        pic[ 715 ] <= 8'd 0 ;
        pic[ 716 ] <= 8'd 0 ;
        pic[ 717 ] <= 8'd 0 ;
        pic[ 718 ] <= 8'd 0 ;
        pic[ 719 ] <= 8'd 0 ;
        pic[ 720 ] <= 8'd 0 ;
        pic[ 721 ] <= 8'd 0 ;
        pic[ 722 ] <= 8'd 0 ;
        pic[ 723 ] <= 8'd 0 ;
        pic[ 724 ] <= 8'd 0 ;
        pic[ 725 ] <= 8'd 0 ;
        pic[ 726 ] <= 8'd 0 ;
        pic[ 727 ] <= 8'd 0 ;
        pic[ 728 ] <= 8'd 0 ;
        pic[ 729 ] <= 8'd 0 ;
        pic[ 730 ] <= 8'd 0 ;
        pic[ 731 ] <= 8'd 0 ;
        pic[ 732 ] <= 8'd 0 ;
        pic[ 733 ] <= 8'd 0 ;
        pic[ 734 ] <= 8'd 0 ;
        pic[ 735 ] <= 8'd 0 ;
        pic[ 736 ] <= 8'd 0 ;
        pic[ 737 ] <= 8'd 0 ;
        pic[ 738 ] <= 8'd 0 ;
        pic[ 739 ] <= 8'd 0 ;
        pic[ 740 ] <= 8'd 0 ;
        pic[ 741 ] <= 8'd 0 ;
        pic[ 742 ] <= 8'd 0 ;
        pic[ 743 ] <= 8'd 0 ;
        pic[ 744 ] <= 8'd 0 ;
        pic[ 745 ] <= 8'd 0 ;
        pic[ 746 ] <= 8'd 0 ;
        pic[ 747 ] <= 8'd 0 ;
        pic[ 748 ] <= 8'd 0 ;
        pic[ 749 ] <= 8'd 0 ;
        pic[ 750 ] <= 8'd 0 ;
        pic[ 751 ] <= 8'd 0 ;
        pic[ 752 ] <= 8'd 0 ;
        pic[ 753 ] <= 8'd 0 ;
        pic[ 754 ] <= 8'd 0 ;
        pic[ 755 ] <= 8'd 0 ;
        pic[ 756 ] <= 8'd 0 ;
        pic[ 757 ] <= 8'd 0 ;
        pic[ 758 ] <= 8'd 0 ;
        pic[ 759 ] <= 8'd 0 ;
        pic[ 760 ] <= 8'd 0 ;
        pic[ 761 ] <= 8'd 0 ;
        pic[ 762 ] <= 8'd 0 ;
        pic[ 763 ] <= 8'd 0 ;
        pic[ 764 ] <= 8'd 0 ;
        pic[ 765 ] <= 8'd 0 ;
        pic[ 766 ] <= 8'd 0 ;
        pic[ 767 ] <= 8'd 0 ;
        pic[ 768 ] <= 8'd 0 ;
        pic[ 769 ] <= 8'd 0 ;
        pic[ 770 ] <= 8'd 0 ;
        pic[ 771 ] <= 8'd 0 ;
        pic[ 772 ] <= 8'd 0 ;
        pic[ 773 ] <= 8'd 0 ;
        pic[ 774 ] <= 8'd 0 ;
        pic[ 775 ] <= 8'd 0 ;
        pic[ 776 ] <= 8'd 0 ;
        pic[ 777 ] <= 8'd 0 ;
        pic[ 778 ] <= 8'd 0 ;
        pic[ 779 ] <= 8'd 0 ;
        pic[ 780 ] <= 8'd 0 ;
        pic[ 781 ] <= 8'd 0 ;
        pic[ 782 ] <= 8'd 0 ;
        pic[ 783 ] <= 8'd 0 ;
		end
		else begin
			for (cnt = 10'd0; cnt < 10'd783; cnt = cnt + 1'd1) begin
				pic[cnt] <= pic[cnt];
			end
			if (addr <= 10'd783)
				data_out <= pic[addr];
			else// invalid addr
				data_out <= 8'd0;
		end
	end
endmodule
