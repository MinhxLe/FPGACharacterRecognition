`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:51:07 05/28/2016 
// Design Name: 
// Module Name:    pic_ram 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module weight_ram(
	clk,
	rst,
	addr,
	data_out
    );
	input clk;
	input rst;
	input [9:0] addr;
	output reg [31:0] data_out;
	reg cnt;
	
	reg [31:0] weights [0:784];

	always @ (posedge clk) begin
		if (rst) begin
			//weights
		  //addr <= 10'd0;
        weights[ 0 ] <= 32'h 38755540 ;
        weights[ 1 ] <= 32'h 0 ;
        weights[ 2 ] <= 32'h 0 ;
        weights[ 3 ] <= 32'h 0 ;
        weights[ 4 ] <= 32'h 0 ;
        weights[ 5 ] <= 32'h 0 ;
        weights[ 6 ] <= 32'h 0 ;
        weights[ 7 ] <= 32'h 0 ;
        weights[ 8 ] <= 32'h 0 ;
        weights[ 9 ] <= 32'h 0 ;
        weights[ 10 ] <= 32'h 0 ;
        weights[ 11 ] <= 32'h 0 ;
        weights[ 12 ] <= 32'h 0 ;
        weights[ 13 ] <= 32'h 0 ;
        weights[ 14 ] <= 32'h 0 ;
        weights[ 15 ] <= 32'h 0 ;
        weights[ 16 ] <= 32'h 0 ;
        weights[ 17 ] <= 32'h 0 ;
        weights[ 18 ] <= 32'h 0 ;
        weights[ 19 ] <= 32'h 0 ;
        weights[ 20 ] <= 32'h 0 ;
        weights[ 21 ] <= 32'h 0 ;
        weights[ 22 ] <= 32'h 0 ;
        weights[ 23 ] <= 32'h 0 ;
        weights[ 24 ] <= 32'h 0 ;
        weights[ 25 ] <= 32'h 0 ;
        weights[ 26 ] <= 32'h 0 ;
        weights[ 27 ] <= 32'h 0 ;
        weights[ 28 ] <= 32'h 0 ;
        weights[ 29 ] <= 32'h 0 ;
        weights[ 30 ] <= 32'h 0 ;
        weights[ 31 ] <= 32'h 0 ;
        weights[ 32 ] <= 32'h 0 ;
        weights[ 33 ] <= 32'h 0 ;
        weights[ 34 ] <= 32'h 0 ;
        weights[ 35 ] <= 32'h 0 ;
        weights[ 36 ] <= 32'h 0 ;
        weights[ 37 ] <= 32'h 0 ;
        weights[ 38 ] <= 32'h 0 ;
        weights[ 39 ] <= 32'h 0 ;
        weights[ 40 ] <= 32'h b628b925 ;
        weights[ 41 ] <= 32'h b6a6befa ;
        weights[ 42 ] <= 32'h b609166e ;
        weights[ 43 ] <= 32'h 36cda1a5 ;
        weights[ 44 ] <= 32'h b9af4c0f ;
        weights[ 45 ] <= 32'h ba765b51 ;
        weights[ 46 ] <= 32'h b9eaafe3 ;
        weights[ 47 ] <= 32'h 0 ;
        weights[ 48 ] <= 32'h 0 ;
        weights[ 49 ] <= 32'h 0 ;
        weights[ 50 ] <= 32'h 0 ;
        weights[ 51 ] <= 32'h 0 ;
        weights[ 52 ] <= 32'h 0 ;
        weights[ 53 ] <= 32'h 0 ;
        weights[ 54 ] <= 32'h 0 ;
        weights[ 55 ] <= 32'h 0 ;
        weights[ 56 ] <= 32'h 0 ;
        weights[ 57 ] <= 32'h 0 ;
        weights[ 58 ] <= 32'h 0 ;
        weights[ 59 ] <= 32'h 0 ;
        weights[ 60 ] <= 32'h b518e7ca ;
        weights[ 61 ] <= 32'h b452e76e ;
        weights[ 62 ] <= 32'h 0 ;
        weights[ 63 ] <= 32'h b5e015e5 ;
        weights[ 64 ] <= 32'h b683d0a5 ;
        weights[ 65 ] <= 32'h b567fe93 ;
        weights[ 66 ] <= 32'h 0 ;
        weights[ 67 ] <= 32'h 35e2b8ca ;
        weights[ 68 ] <= 32'h 3771df66 ;
        weights[ 69 ] <= 32'h 3987db71 ;
        weights[ 70 ] <= 32'h 3ab229eb ;
        weights[ 71 ] <= 32'h 3a7bb457 ;
        weights[ 72 ] <= 32'h 3a5c7d80 ;
        weights[ 73 ] <= 32'h 3a15f192 ;
        weights[ 74 ] <= 32'h 3a7a0dae ;
        weights[ 75 ] <= 32'h 3986a19e ;
        weights[ 76 ] <= 32'h 38963e1f ;
        weights[ 77 ] <= 32'h 3793d643 ;
        weights[ 78 ] <= 32'h 0 ;
        weights[ 79 ] <= 32'h 0 ;
        weights[ 80 ] <= 32'h 0 ;
        weights[ 81 ] <= 32'h 0 ;
        weights[ 82 ] <= 32'h 0 ;
        weights[ 83 ] <= 32'h 0 ;
        weights[ 84 ] <= 32'h 0 ;
        weights[ 85 ] <= 32'h 0 ;
        weights[ 86 ] <= 32'h 0 ;
        weights[ 87 ] <= 32'h 355d7301 ;
        weights[ 88 ] <= 32'h b5c31613 ;
        weights[ 89 ] <= 32'h b623735c ;
        weights[ 90 ] <= 32'h b6ff0fe3 ;
        weights[ 91 ] <= 32'h b6da2763 ;
        weights[ 92 ] <= 32'h b6dec473 ;
        weights[ 93 ] <= 32'h 386fd095 ;
        weights[ 94 ] <= 32'h 39046071 ;
        weights[ 95 ] <= 32'h 385d5ec9 ;
        weights[ 96 ] <= 32'h 393135c4 ;
        weights[ 97 ] <= 32'h 3a91fe04 ;
        weights[ 98 ] <= 32'h 3b20ca5a ;
        weights[ 99 ] <= 32'h 3b846a0d ;
        weights[ 100 ] <= 32'h 3b3f151d ;
        weights[ 101 ] <= 32'h 3b34ebb6 ;
        weights[ 102 ] <= 32'h 3affc79b ;
        weights[ 103 ] <= 32'h 3a3506a6 ;
        weights[ 104 ] <= 32'h 39ddbf83 ;
        weights[ 105 ] <= 32'h 3a0a1763 ;
        weights[ 106 ] <= 32'h 398fb6e7 ;
        weights[ 107 ] <= 32'h b7b24795 ;
        weights[ 108 ] <= 32'h b738dedd ;
        weights[ 109 ] <= 32'h b6a8106c ;
        weights[ 110 ] <= 32'h b5c0732e ;
        weights[ 111 ] <= 32'h 0 ;
        weights[ 112 ] <= 32'h 0 ;
        weights[ 113 ] <= 32'h 0 ;
        weights[ 114 ] <= 32'h 0 ;
        weights[ 115 ] <= 32'h 363dd04a ;
        weights[ 116 ] <= 32'h b6261640 ;
        weights[ 117 ] <= 32'h 36b929c6 ;
        weights[ 118 ] <= 32'h 38bf7485 ;
        weights[ 119 ] <= 32'h 384dae37 ;
        weights[ 120 ] <= 32'h 3801dbb7 ;
        weights[ 121 ] <= 32'h 3a3c5a74 ;
        weights[ 122 ] <= 32'h 3a9b45d1 ;
        weights[ 123 ] <= 32'h 3a6b13cf ;
        weights[ 124 ] <= 32'h 3a8df1b3 ;
        weights[ 125 ] <= 32'h 3b03f193 ;
        weights[ 126 ] <= 32'h 3b677879 ;
        weights[ 127 ] <= 32'h 3b98662b ;
        weights[ 128 ] <= 32'h 3b644813 ;
        weights[ 129 ] <= 32'h 3a9cfa15 ;
        weights[ 130 ] <= 32'h b9da17d9 ;
        weights[ 131 ] <= 32'h bb042eb7 ;
        weights[ 132 ] <= 32'h 39f1ec5f ;
        weights[ 133 ] <= 32'h 3b1d79e0 ;
        weights[ 134 ] <= 32'h 3aecc038 ;
        weights[ 135 ] <= 32'h 3a28bb1e ;
        weights[ 136 ] <= 32'h 39b08fac ;
        weights[ 137 ] <= 32'h 3821ee50 ;
        weights[ 138 ] <= 32'h b6640a3c ;
        weights[ 139 ] <= 32'h 0 ;
        weights[ 140 ] <= 32'h 0 ;
        weights[ 141 ] <= 32'h 0 ;
        weights[ 142 ] <= 32'h 0 ;
        weights[ 143 ] <= 32'h 35fd15b8 ;
        weights[ 144 ] <= 32'h b509166e ;
        weights[ 145 ] <= 32'h 379447fe ;
        weights[ 146 ] <= 32'h 398f4f75 ;
        weights[ 147 ] <= 32'h 398fc8f5 ;
        weights[ 148 ] <= 32'h 397393b0 ;
        weights[ 149 ] <= 32'h 3a9a6031 ;
        weights[ 150 ] <= 32'h 3b0a5eeb ;
        weights[ 151 ] <= 32'h 3a6d94a4 ;
        weights[ 152 ] <= 32'h b8d38d29 ;
        weights[ 153 ] <= 32'h 3a0db797 ;
        weights[ 154 ] <= 32'h 3b1de313 ;
        weights[ 155 ] <= 32'h 3ad19472 ;
        weights[ 156 ] <= 32'h ba999425 ;
        weights[ 157 ] <= 32'h bb7386a6 ;
        weights[ 158 ] <= 32'h bbb32d17 ;
        weights[ 159 ] <= 32'h bbb2d2b0 ;
        weights[ 160 ] <= 32'h bb0103f9 ;
        weights[ 161 ] <= 32'h 3ae63c13 ;
        weights[ 162 ] <= 32'h 3b25a941 ;
        weights[ 163 ] <= 32'h 3ab5c9d5 ;
        weights[ 164 ] <= 32'h 3af08224 ;
        weights[ 165 ] <= 32'h 3a846f09 ;
        weights[ 166 ] <= 32'h b5d8175f ;
        weights[ 167 ] <= 32'h 358bb953 ;
        weights[ 168 ] <= 32'h 0 ;
        weights[ 169 ] <= 32'h 0 ;
        weights[ 170 ] <= 32'h 0 ;
        weights[ 171 ] <= 32'h 34c85bdc ;
        weights[ 172 ] <= 32'h 36db78d5 ;
        weights[ 173 ] <= 32'h b591cc6e ;
        weights[ 174 ] <= 32'h 390542d4 ;
        weights[ 175 ] <= 32'h 3a15e1b6 ;
        weights[ 176 ] <= 32'h 3aaf64a7 ;
        weights[ 177 ] <= 32'h 3aa17f9d ;
        weights[ 178 ] <= 32'h b89f8c7f ;
        weights[ 179 ] <= 32'h baffdd7d ;
        weights[ 180 ] <= 32'h bb8362e7 ;
        weights[ 181 ] <= 32'h bb4d03fc ;
        weights[ 182 ] <= 32'h bb0fb6ce ;
        weights[ 183 ] <= 32'h bb39d4ff ;
        weights[ 184 ] <= 32'h bb8c3499 ;
        weights[ 185 ] <= 32'h bbe865da ;
        weights[ 186 ] <= 32'h bc08b350 ;
        weights[ 187 ] <= 32'h bbe6174b ;
        weights[ 188 ] <= 32'h bbae76db ;
        weights[ 189 ] <= 32'h bae3bce8 ;
        weights[ 190 ] <= 32'h ba36a95a ;
        weights[ 191 ] <= 32'h ba7480fa ;
        weights[ 192 ] <= 32'h 39c24428 ;
        weights[ 193 ] <= 32'h 3aa91a95 ;
        weights[ 194 ] <= 32'h b6fbc445 ;
        weights[ 195 ] <= 32'h b5d82d37 ;
        weights[ 196 ] <= 32'h b5c0732e ;
        weights[ 197 ] <= 32'h 0 ;
        weights[ 198 ] <= 32'h 0 ;
        weights[ 199 ] <= 32'h 35bdd04a ;
        weights[ 200 ] <= 32'h 352dfeee ;
        weights[ 201 ] <= 32'h 3a28dd57 ;
        weights[ 202 ] <= 32'h 3a4100d4 ;
        weights[ 203 ] <= 32'h 3a86288c ;
        weights[ 204 ] <= 32'h 3b20eeb0 ;
        weights[ 205 ] <= 32'h 398730e7 ;
        weights[ 206 ] <= 32'h bb5269fa ;
        weights[ 207 ] <= 32'h bbd5daea ;
        weights[ 208 ] <= 32'h bc0629c4 ;
        weights[ 209 ] <= 32'h bbd25572 ;
        weights[ 210 ] <= 32'h bb8d587e ;
        weights[ 211 ] <= 32'h bb80a741 ;
        weights[ 212 ] <= 32'h bb3ee69d ;
        weights[ 213 ] <= 32'h bbb1598d ;
        weights[ 214 ] <= 32'h bbfd6bec ;
        weights[ 215 ] <= 32'h bbf1ce8a ;
        weights[ 216 ] <= 32'h bc0a9782 ;
        weights[ 217 ] <= 32'h bbe2f694 ;
        weights[ 218 ] <= 32'h bbc395c4 ;
        weights[ 219 ] <= 32'h bb89f211 ;
        weights[ 220 ] <= 32'h baca831d ;
        weights[ 221 ] <= 32'h 35f0a212 ;
        weights[ 222 ] <= 32'h b7a0a649 ;
        weights[ 223 ] <= 32'h 34e7fe93 ;
        weights[ 224 ] <= 32'h b64afec1 ;
        weights[ 225 ] <= 32'h b58bb953 ;
        weights[ 226 ] <= 32'h 0 ;
        weights[ 227 ] <= 32'h b5c5b8f7 ;
        weights[ 228 ] <= 32'h b577cfee ;
        weights[ 229 ] <= 32'h 3a1d38d0 ;
        weights[ 230 ] <= 32'h 3a43cef8 ;
        weights[ 231 ] <= 32'h 3a7fa36c ;
        weights[ 232 ] <= 32'h 3af29fd2 ;
        weights[ 233 ] <= 32'h b9b79062 ;
        weights[ 234 ] <= 32'h bba28202 ;
        weights[ 235 ] <= 32'h bbf80837 ;
        weights[ 236 ] <= 32'h bbffda43 ;
        weights[ 237 ] <= 32'h bbc812a6 ;
        weights[ 238 ] <= 32'h bb9d2561 ;
        weights[ 239 ] <= 32'h 38c0aa58 ;
        weights[ 240 ] <= 32'h 3b48f307 ;
        weights[ 241 ] <= 32'h ba4c04b3 ;
        weights[ 242 ] <= 32'h bb9f0097 ;
        weights[ 243 ] <= 32'h bbfa51a8 ;
        weights[ 244 ] <= 32'h bc2a746b ;
        weights[ 245 ] <= 32'h bc40c109 ;
        weights[ 246 ] <= 32'h bc37ace8 ;
        weights[ 247 ] <= 32'h bbf7ee38 ;
        weights[ 248 ] <= 32'h bb5382e1 ;
        weights[ 249 ] <= 32'h ba273b72 ;
        weights[ 250 ] <= 32'h b773db98 ;
        weights[ 251 ] <= 32'h 0 ;
        weights[ 252 ] <= 32'h 0 ;
        weights[ 253 ] <= 32'h 0 ;
        weights[ 254 ] <= 32'h 35d58a53 ;
        weights[ 255 ] <= 32'h b562b8ca ;
        weights[ 256 ] <= 32'h b69cdc20 ;
        weights[ 257 ] <= 32'h 3a3cd8c3 ;
        weights[ 258 ] <= 32'h 39ffec9d ;
        weights[ 259 ] <= 32'h b9d5a79f ;
        weights[ 260 ] <= 32'h 39a23ef4 ;
        weights[ 261 ] <= 32'h badfeb20 ;
        weights[ 262 ] <= 32'h bba1af7c ;
        weights[ 263 ] <= 32'h bbed451e ;
        weights[ 264 ] <= 32'h bbfaf259 ;
        weights[ 265 ] <= 32'h bbdd0b88 ;
        weights[ 266 ] <= 32'h bb138fe1 ;
        weights[ 267 ] <= 32'h 3bc20503 ;
        weights[ 268 ] <= 32'h 3c306edc ;
        weights[ 269 ] <= 32'h 3bf19b32 ;
        weights[ 270 ] <= 32'h 3a6bac06 ;
        weights[ 271 ] <= 32'h bb984ea1 ;
        weights[ 272 ] <= 32'h bc1f7b51 ;
        weights[ 273 ] <= 32'h bc70f5c3 ;
        weights[ 274 ] <= 32'h bc8162dd ;
        weights[ 275 ] <= 32'h bc348461 ;
        weights[ 276 ] <= 32'h bbb5627f ;
        weights[ 277 ] <= 32'h baae3cb1 ;
        weights[ 278 ] <= 32'h b78994f9 ;
        weights[ 279 ] <= 32'h 35a61640 ;
        weights[ 280 ] <= 32'h 0 ;
        weights[ 281 ] <= 32'h 0 ;
        weights[ 282 ] <= 32'h 362f5061 ;
        weights[ 283 ] <= 32'h b637390e ;
        weights[ 284 ] <= 32'h b69cdc20 ;
        weights[ 285 ] <= 32'h 3a32c676 ;
        weights[ 286 ] <= 32'h b99b196a ;
        weights[ 287 ] <= 32'h bacc8a47 ;
        weights[ 288 ] <= 32'h bb5f9301 ;
        weights[ 289 ] <= 32'h bbb03543 ;
        weights[ 290 ] <= 32'h bbe87886 ;
        weights[ 291 ] <= 32'h bc0b8216 ;
        weights[ 292 ] <= 32'h bc1301e2 ;
        weights[ 293 ] <= 32'h bc024a44 ;
        weights[ 294 ] <= 32'h ba29caa8 ;
        weights[ 295 ] <= 32'h 3c3fba34 ;
        weights[ 296 ] <= 32'h 3c9c5c1e ;
        weights[ 297 ] <= 32'h 3c4ce7a3 ;
        weights[ 298 ] <= 32'h 3b8cc72f ;
        weights[ 299 ] <= 32'h bb133a73 ;
        weights[ 300 ] <= 32'h bc1b11c1 ;
        weights[ 301 ] <= 32'h bc8c9cf1 ;
        weights[ 302 ] <= 32'h bc913c8e ;
        weights[ 303 ] <= 32'h bc5f1b44 ;
        weights[ 304 ] <= 32'h bbf1aa57 ;
        weights[ 305 ] <= 32'h bb02896d ;
        weights[ 306 ] <= 32'h b7f72735 ;
        weights[ 307 ] <= 32'h 36640a3c ;
        weights[ 308 ] <= 32'h 35485bdc ;
        weights[ 309 ] <= 32'h 0 ;
        weights[ 310 ] <= 32'h 3518e7ca ;
        weights[ 311 ] <= 32'h 35485bdc ;
        weights[ 312 ] <= 32'h b637390e ;
        weights[ 313 ] <= 32'h 3a1bb131 ;
        weights[ 314 ] <= 32'h ba736f24 ;
        weights[ 315 ] <= 32'h bb4fafd8 ;
        weights[ 316 ] <= 32'h bbd8495c ;
        weights[ 317 ] <= 32'h bc218184 ;
        weights[ 318 ] <= 32'h bc37b876 ;
        weights[ 319 ] <= 32'h bc4066ea ;
        weights[ 320 ] <= 32'h bc44c8b7 ;
        weights[ 321 ] <= 32'h bc0c951c ;
        weights[ 322 ] <= 32'h 3b54c034 ;
        weights[ 323 ] <= 32'h 3ca0c6cf ;
        weights[ 324 ] <= 32'h 3cd14f08 ;
        weights[ 325 ] <= 32'h 3c8a17b7 ;
        weights[ 326 ] <= 32'h 3babd410 ;
        weights[ 327 ] <= 32'h bb35e84f ;
        weights[ 328 ] <= 32'h bc3288fb ;
        weights[ 329 ] <= 32'h bc867048 ;
        weights[ 330 ] <= 32'h bc91ca16 ;
        weights[ 331 ] <= 32'h bc6e8029 ;
        weights[ 332 ] <= 32'h bc09fa40 ;
        weights[ 333 ] <= 32'h bb2ee001 ;
        weights[ 334 ] <= 32'h b86c322f ;
        weights[ 335 ] <= 32'h b5a61640 ;
        weights[ 336 ] <= 32'h 35efe741 ;
        weights[ 337 ] <= 32'h 0 ;
        weights[ 338 ] <= 32'h b4a8b925 ;
        weights[ 339 ] <= 32'h b57d15b8 ;
        weights[ 340 ] <= 32'h b3fd15b8 ;
        weights[ 341 ] <= 32'h 39cd32c4 ;
        weights[ 342 ] <= 32'h bb121ac3 ;
        weights[ 343 ] <= 32'h bbada448 ;
        weights[ 344 ] <= 32'h bc1b1684 ;
        weights[ 345 ] <= 32'h bc5742a8 ;
        weights[ 346 ] <= 32'h bc6961a9 ;
        weights[ 347 ] <= 32'h bc65c64f ;
        weights[ 348 ] <= 32'h bc461f9f ;
        weights[ 349 ] <= 32'h bc0e9c8b ;
        weights[ 350 ] <= 32'h 3c09b24c ;
        weights[ 351 ] <= 32'h 3ce48655 ;
        weights[ 352 ] <= 32'h 3cf85ca3 ;
        weights[ 353 ] <= 32'h 3c96bd61 ;
        weights[ 354 ] <= 32'h 3b82c7d4 ;
        weights[ 355 ] <= 32'h bb9fa7a0 ;
        weights[ 356 ] <= 32'h bc3ecd54 ;
        weights[ 357 ] <= 32'h bc81942c ;
        weights[ 358 ] <= 32'h bc90d804 ;
        weights[ 359 ] <= 32'h bc787209 ;
        weights[ 360 ] <= 32'h bc1f4b67 ;
        weights[ 361 ] <= 32'h bb562098 ;
        weights[ 362 ] <= 32'h b8b8bf3a ;
        weights[ 363 ] <= 32'h b64c5033 ;
        weights[ 364 ] <= 32'h 3610ff1c ;
        weights[ 365 ] <= 32'h 3528b925 ;
        weights[ 366 ] <= 32'h b5a61640 ;
        weights[ 367 ] <= 32'h b65c218e ;
        weights[ 368 ] <= 32'h b6d438e1 ;
        weights[ 369 ] <= 32'h b9a95a1a ;
        weights[ 370 ] <= 32'h bb76e602 ;
        weights[ 371 ] <= 32'h bc02c7d0 ;
        weights[ 372 ] <= 32'h bc5876f6 ;
        weights[ 373 ] <= 32'h bc88b377 ;
        weights[ 374 ] <= 32'h bc900f1a ;
        weights[ 375 ] <= 32'h bc710eb0 ;
        weights[ 376 ] <= 32'h bc4c85bd ;
        weights[ 377 ] <= 32'h bbd44d0c ;
        weights[ 378 ] <= 32'h 3c86ecec ;
        weights[ 379 ] <= 32'h 3d07f9bd ;
        weights[ 380 ] <= 32'h 3d04d1b3 ;
        weights[ 381 ] <= 32'h 3c899dfb ;
        weights[ 382 ] <= 32'h 3b09a9f7 ;
        weights[ 383 ] <= 32'h bc040481 ;
        weights[ 384 ] <= 32'h bc4900aa ;
        weights[ 385 ] <= 32'h bc7cbcb9 ;
        weights[ 386 ] <= 32'h bc9545d0 ;
        weights[ 387 ] <= 32'h bc821cfa ;
        weights[ 388 ] <= 32'h bc28947c ;
        weights[ 389 ] <= 32'h bb6ae8fa ;
        weights[ 390 ] <= 32'h b9000137 ;
        weights[ 391 ] <= 32'h b3fd15b8 ;
        weights[ 392 ] <= 32'h 0 ;
        weights[ 393 ] <= 32'h 0 ;
        weights[ 394 ] <= 32'h 0 ;
        weights[ 395 ] <= 32'h 3467fe93 ;
        weights[ 396 ] <= 32'h b53dd04a ;
        weights[ 397 ] <= 32'h ba33d9c5 ;
        weights[ 398 ] <= 32'h bbb188e7 ;
        weights[ 399 ] <= 32'h bc3e3b22 ;
        weights[ 400 ] <= 32'h bc8d09cd ;
        weights[ 401 ] <= 32'h bc986361 ;
        weights[ 402 ] <= 32'h bc80d7d4 ;
        weights[ 403 ] <= 32'h bc6e2ab2 ;
        weights[ 404 ] <= 32'h bc36b7d7 ;
        weights[ 405 ] <= 32'h b9b1668b ;
        weights[ 406 ] <= 32'h 3cbd1339 ;
        weights[ 407 ] <= 32'h 3d147971 ;
        weights[ 408 ] <= 32'h 3d023eb2 ;
        weights[ 409 ] <= 32'h 3c4fcc5f ;
        weights[ 410 ] <= 32'h ba7d595c ;
        weights[ 411 ] <= 32'h bc21b188 ;
        weights[ 412 ] <= 32'h bc4ec517 ;
        weights[ 413 ] <= 32'h bc8200d9 ;
        weights[ 414 ] <= 32'h bc93e4d1 ;
        weights[ 415 ] <= 32'h bc791978 ;
        weights[ 416 ] <= 32'h bc1fb662 ;
        weights[ 417 ] <= 32'h bb694db7 ;
        weights[ 418 ] <= 32'h b91970e0 ;
        weights[ 419 ] <= 32'h 3503d0a5 ;
        weights[ 420 ] <= 32'h 0 ;
        weights[ 421 ] <= 32'h 0 ;
        weights[ 422 ] <= 32'h 0 ;
        weights[ 423 ] <= 32'h 35fa72d3 ;
        weights[ 424 ] <= 32'h b66d445c ;
        weights[ 425 ] <= 32'h bacd9e5a ;
        weights[ 426 ] <= 32'h bbfb6e6d ;
        weights[ 427 ] <= 32'h bc676dfd ;
        weights[ 428 ] <= 32'h bc985d30 ;
        weights[ 429 ] <= 32'h bc93a8a5 ;
        weights[ 430 ] <= 32'h bc7e3955 ;
        weights[ 431 ] <= 32'h bc6ad288 ;
        weights[ 432 ] <= 32'h bbfce3c8 ;
        weights[ 433 ] <= 32'h 3bf5db79 ;
        weights[ 434 ] <= 32'h 3ce0614c ;
        weights[ 435 ] <= 32'h 3d1896bf ;
        weights[ 436 ] <= 32'h 3cdd75bf ;
        weights[ 437 ] <= 32'h 3bf640f4 ;
        weights[ 438 ] <= 32'h bb96f4e8 ;
        weights[ 439 ] <= 32'h bc1d3930 ;
        weights[ 440 ] <= 32'h bc5e1f70 ;
        weights[ 441 ] <= 32'h bc84a7f2 ;
        weights[ 442 ] <= 32'h bc8d7b1e ;
        weights[ 443 ] <= 32'h bc65ba03 ;
        weights[ 444 ] <= 32'h bc0cfe7f ;
        weights[ 445 ] <= 32'h bb488119 ;
        weights[ 446 ] <= 32'h b9074bb7 ;
        weights[ 447 ] <= 32'h 3452e76e ;
        weights[ 448 ] <= 32'h 0 ;
        weights[ 449 ] <= 32'h 0 ;
        weights[ 450 ] <= 32'h 354da1a5 ;
        weights[ 451 ] <= 32'h 3645b8f7 ;
        weights[ 452 ] <= 32'h b7777b92 ;
        weights[ 453 ] <= 32'h bb0d9fb8 ;
        weights[ 454 ] <= 32'h bc167bc3 ;
        weights[ 455 ] <= 32'h bc801987 ;
        weights[ 456 ] <= 32'h bc9d6164 ;
        weights[ 457 ] <= 32'h bc911efc ;
        weights[ 458 ] <= 32'h bc83b1a9 ;
        weights[ 459 ] <= 32'h bc3dc41f ;
        weights[ 460 ] <= 32'h bb058cc7 ;
        weights[ 461 ] <= 32'h 3c52f125 ;
        weights[ 462 ] <= 32'h 3ce79184 ;
        weights[ 463 ] <= 32'h 3d046b6a ;
        weights[ 464 ] <= 32'h 3ca7583c ;
        weights[ 465 ] <= 32'h 3b33fcdc ;
        weights[ 466 ] <= 32'h bbdbe185 ;
        weights[ 467 ] <= 32'h bc1dba66 ;
        weights[ 468 ] <= 32'h bc646a26 ;
        weights[ 469 ] <= 32'h bc885fc7 ;
        weights[ 470 ] <= 32'h bc80cc10 ;
        weights[ 471 ] <= 32'h bc4280b7 ;
        weights[ 472 ] <= 32'h bbd89215 ;
        weights[ 473 ] <= 32'h bac88719 ;
        weights[ 474 ] <= 32'h 3918ee5b ;
        weights[ 475 ] <= 32'h 3640732e ;
        weights[ 476 ] <= 32'h b47d15b8 ;
        weights[ 477 ] <= 32'h 0 ;
        weights[ 478 ] <= 32'h 362767b3 ;
        weights[ 479 ] <= 32'h 3567fe93 ;
        weights[ 480 ] <= 32'h b7d29312 ;
        weights[ 481 ] <= 32'h bb34f85d ;
        weights[ 482 ] <= 32'h bc259e77 ;
        weights[ 483 ] <= 32'h bc83c694 ;
        weights[ 484 ] <= 32'h bc93f54f ;
        weights[ 485 ] <= 32'h bc8e2023 ;
        weights[ 486 ] <= 32'h bc72051c ;
        weights[ 487 ] <= 32'h bc01aa26 ;
        weights[ 488 ] <= 32'h 3b15f1ee ;
        weights[ 489 ] <= 32'h 3c759ebb ;
        weights[ 490 ] <= 32'h 3cd074fa ;
        weights[ 491 ] <= 32'h 3cd0867a ;
        weights[ 492 ] <= 32'h 3c6f1fb1 ;
        weights[ 493 ] <= 32'h b8d26760 ;
        weights[ 494 ] <= 32'h bc0e8d19 ;
        weights[ 495 ] <= 32'h bc35d9c8 ;
        weights[ 496 ] <= 32'h bc6af045 ;
        weights[ 497 ] <= 32'h bc82a820 ;
        weights[ 498 ] <= 32'h bc532473 ;
        weights[ 499 ] <= 32'h bc0d05f8 ;
        weights[ 500 ] <= 32'h bb8ad7c6 ;
        weights[ 501 ] <= 32'h b98797ad ;
        weights[ 502 ] <= 32'h 3a77e5c0 ;
        weights[ 503 ] <= 32'h 369d84da ;
        weights[ 504 ] <= 32'h b5fd15b8 ;
        weights[ 505 ] <= 32'h 337d15b8 ;
        weights[ 506 ] <= 32'h 34fd15b8 ;
        weights[ 507 ] <= 32'h 33d2e76e ;
        weights[ 508 ] <= 32'h b812f947 ;
        weights[ 509 ] <= 32'h bb45308a ;
        weights[ 510 ] <= 32'h bc23cf30 ;
        weights[ 511 ] <= 32'h bc794d6a ;
        weights[ 512 ] <= 32'h bc8df936 ;
        weights[ 513 ] <= 32'h bc9182fc ;
        weights[ 514 ] <= 32'h bc607df7 ;
        weights[ 515 ] <= 32'h bbba73e3 ;
        weights[ 516 ] <= 32'h 3b4e3367 ;
        weights[ 517 ] <= 32'h 3c66122f ;
        weights[ 518 ] <= 32'h 3cafb25c ;
        weights[ 519 ] <= 32'h 3c91fcf1 ;
        weights[ 520 ] <= 32'h 3beeda0a ;
        weights[ 521 ] <= 32'h bb538f38 ;
        weights[ 522 ] <= 32'h bc238ee2 ;
        weights[ 523 ] <= 32'h bc406fce ;
        weights[ 524 ] <= 32'h bc67bc3b ;
        weights[ 525 ] <= 32'h bc491d19 ;
        weights[ 526 ] <= 32'h bc118581 ;
        weights[ 527 ] <= 32'h bbae0f28 ;
        weights[ 528 ] <= 32'h bac824cb ;
        weights[ 529 ] <= 32'h 3a69241a ;
        weights[ 530 ] <= 32'h 3a86fda9 ;
        weights[ 531 ] <= 32'h 36e2b8ca ;
        weights[ 532 ] <= 32'h 369ed64c ;
        weights[ 533 ] <= 32'h 349e2d93 ;
        weights[ 534 ] <= 32'h 351e2c17 ;
        weights[ 535 ] <= 32'h b4891956 ;
        weights[ 536 ] <= 32'h b840b278 ;
        weights[ 537 ] <= 32'h bb37d73c ;
        weights[ 538 ] <= 32'h bc114261 ;
        weights[ 539 ] <= 32'h bc54f018 ;
        weights[ 540 ] <= 32'h bc7f18f1 ;
        weights[ 541 ] <= 32'h bc857bb7 ;
        weights[ 542 ] <= 32'h bc46e892 ;
        weights[ 543 ] <= 32'h bb81c67e ;
        weights[ 544 ] <= 32'h 3b7d1c7a ;
        weights[ 545 ] <= 32'h 3c3e9fce ;
        weights[ 546 ] <= 32'h 3c8089d2 ;
        weights[ 547 ] <= 32'h 3c3c50c6 ;
        weights[ 548 ] <= 32'h 3b354ff3 ;
        weights[ 549 ] <= 32'h bb8668df ;
        weights[ 550 ] <= 32'h bc08e8b0 ;
        weights[ 551 ] <= 32'h bc220c78 ;
        weights[ 552 ] <= 32'h bc19de51 ;
        weights[ 553 ] <= 32'h bbdc4ff0 ;
        weights[ 554 ] <= 32'h bb80afc8 ;
        weights[ 555 ] <= 32'h ba8efb55 ;
        weights[ 556 ] <= 32'h 3a8dc195 ;
        weights[ 557 ] <= 32'h 3afad363 ;
        weights[ 558 ] <= 32'h 3a8a0821 ;
        weights[ 559 ] <= 32'h 368fadaa ;
        weights[ 560 ] <= 32'h 365438e1 ;
        weights[ 561 ] <= 32'h 0 ;
        weights[ 562 ] <= 32'h b62cae6b ;
        weights[ 563 ] <= 32'h b5d82e84 ;
        weights[ 564 ] <= 32'h 38a8df68 ;
        weights[ 565 ] <= 32'h bafd966c ;
        weights[ 566 ] <= 32'h bbc102f9 ;
        weights[ 567 ] <= 32'h bc0b48f2 ;
        weights[ 568 ] <= 32'h bc3d0a28 ;
        weights[ 569 ] <= 32'h bc4afbb3 ;
        weights[ 570 ] <= 32'h bc16a0c5 ;
        weights[ 571 ] <= 32'h bb740600 ;
        weights[ 572 ] <= 32'h 3aeab932 ;
        weights[ 573 ] <= 32'h 3bc7256b ;
        weights[ 574 ] <= 32'h 3bf57616 ;
        weights[ 575 ] <= 32'h 3bbc6e63 ;
        weights[ 576 ] <= 32'h 398501c6 ;
        weights[ 577 ] <= 32'h bb80c60e ;
        weights[ 578 ] <= 32'h bb793ae8 ;
        weights[ 579 ] <= 32'h bb3a0341 ;
        weights[ 580 ] <= 32'h bab66cc5 ;
        weights[ 581 ] <= 32'h 39cdf00c ;
        weights[ 582 ] <= 32'h 3a48e46a ;
        weights[ 583 ] <= 32'h 3b01edbb ;
        weights[ 584 ] <= 32'h 3b33ac5c ;
        weights[ 585 ] <= 32'h 3b1d49c0 ;
        weights[ 586 ] <= 32'h 3a708b0e ;
        weights[ 587 ] <= 32'h 35728a25 ;
        weights[ 588 ] <= 32'h 3586738a ;
        weights[ 589 ] <= 32'h 3528b925 ;
        weights[ 590 ] <= 32'h 3452e76e ;
        weights[ 591 ] <= 32'h 35485bdc ;
        weights[ 592 ] <= 32'h 3a03a4c7 ;
        weights[ 593 ] <= 32'h 3a3e5407 ;
        weights[ 594 ] <= 32'h 3a8ada3a ;
        weights[ 595 ] <= 32'h ba94168f ;
        weights[ 596 ] <= 32'h bb89304e ;
        weights[ 597 ] <= 32'h bbce3235 ;
        weights[ 598 ] <= 32'h bbccd44d ;
        weights[ 599 ] <= 32'h bbad494a ;
        weights[ 600 ] <= 32'h bb70b84f ;
        weights[ 601 ] <= 32'h ba6a5576 ;
        weights[ 602 ] <= 32'h 3ae17466 ;
        weights[ 603 ] <= 32'h 3a7335a6 ;
        weights[ 604 ] <= 32'h bb02b548 ;
        weights[ 605 ] <= 32'h bb12c5dc ;
        weights[ 606 ] <= 32'h ba8117d6 ;
        weights[ 607 ] <= 32'h 3a44cc47 ;
        weights[ 608 ] <= 32'h 3b13ec7c ;
        weights[ 609 ] <= 32'h 3ba0382e ;
        weights[ 610 ] <= 32'h 3b94ee14 ;
        weights[ 611 ] <= 32'h 3b174205 ;
        weights[ 612 ] <= 32'h 3af088a0 ;
        weights[ 613 ] <= 32'h 3b0397c8 ;
        weights[ 614 ] <= 32'h 3a92094e ;
        weights[ 615 ] <= 32'h b68f04f0 ;
        weights[ 616 ] <= 32'h b54da1a5 ;
        weights[ 617 ] <= 32'h 3523735c ;
        weights[ 618 ] <= 32'h 3452e76e ;
        weights[ 619 ] <= 32'h 35c5b8f7 ;
        weights[ 620 ] <= 32'h 3968d405 ;
        weights[ 621 ] <= 32'h 3b097d2e ;
        weights[ 622 ] <= 32'h 3b45f25b ;
        weights[ 623 ] <= 32'h 3ac1d02e ;
        weights[ 624 ] <= 32'h baae63ab ;
        weights[ 625 ] <= 32'h bb2f0dbc ;
        weights[ 626 ] <= 32'h bb7e4979 ;
        weights[ 627 ] <= 32'h bbcf7ed9 ;
        weights[ 628 ] <= 32'h bc0a33c9 ;
        weights[ 629 ] <= 32'h bbf1af4b ;
        weights[ 630 ] <= 32'h bba15ebd ;
        weights[ 631 ] <= 32'h bb6c4a7e ;
        weights[ 632 ] <= 32'h bb5a7608 ;
        weights[ 633 ] <= 32'h bb2d69fa ;
        weights[ 634 ] <= 32'h baf28065 ;
        weights[ 635 ] <= 32'h b8baeae1 ;
        weights[ 636 ] <= 32'h 3a8e2a05 ;
        weights[ 637 ] <= 32'h 3b554025 ;
        weights[ 638 ] <= 32'h 3b448b76 ;
        weights[ 639 ] <= 32'h 3a5609be ;
        weights[ 640 ] <= 32'h 3a08ef19 ;
        weights[ 641 ] <= 32'h 3a1ae0f9 ;
        weights[ 642 ] <= 32'h 3a04c94c ;
        weights[ 643 ] <= 32'h 36012dc0 ;
        weights[ 644 ] <= 32'h b5bdd04a ;
        weights[ 645 ] <= 32'h 0 ;
        weights[ 646 ] <= 32'h 0 ;
        weights[ 647 ] <= 32'h 0 ;
        weights[ 648 ] <= 32'h b577cfee ;
        weights[ 649 ] <= 32'h 39cfc9ac ;
        weights[ 650 ] <= 32'h 3a05ccfb ;
        weights[ 651 ] <= 32'h 3a200492 ;
        weights[ 652 ] <= 32'h ba0e5336 ;
        weights[ 653 ] <= 32'h ba672e26 ;
        weights[ 654 ] <= 32'h ba651dd1 ;
        weights[ 655 ] <= 32'h bba6c6d3 ;
        weights[ 656 ] <= 32'h bc18aabf ;
        weights[ 657 ] <= 32'h bc082c74 ;
        weights[ 658 ] <= 32'h bbae8b7d ;
        weights[ 659 ] <= 32'h bb6e366b ;
        weights[ 660 ] <= 32'h baf6eda2 ;
        weights[ 661 ] <= 32'h bafd8d26 ;
        weights[ 662 ] <= 32'h bb0132b0 ;
        weights[ 663 ] <= 32'h ba6a6672 ;
        weights[ 664 ] <= 32'h 39b403a5 ;
        weights[ 665 ] <= 32'h 3aad473d ;
        weights[ 666 ] <= 32'h 3a0f283b ;
        weights[ 667 ] <= 32'h 38c1cd68 ;
        weights[ 668 ] <= 32'h b71c50aa ;
        weights[ 669 ] <= 32'h b61644e5 ;
        weights[ 670 ] <= 32'h 3650448a ;
        weights[ 671 ] <= 32'h 36bf21bc ;
        weights[ 672 ] <= 32'h 0 ;
        weights[ 673 ] <= 32'h 0 ;
        weights[ 674 ] <= 32'h 0 ;
        weights[ 675 ] <= 32'h 0 ;
        weights[ 676 ] <= 32'h 32a8b925 ;
        weights[ 677 ] <= 32'h b47bd296 ;
        weights[ 678 ] <= 32'h 3902ea23 ;
        weights[ 679 ] <= 32'h 399ac6fb ;
        weights[ 680 ] <= 32'h 3a4da5b6 ;
        weights[ 681 ] <= 32'h 3a456835 ;
        weights[ 682 ] <= 32'h 3a6d30e2 ;
        weights[ 683 ] <= 32'h 39b41a14 ;
        weights[ 684 ] <= 32'h bac33936 ;
        weights[ 685 ] <= 32'h bb3edc3a ;
        weights[ 686 ] <= 32'h bb10218b ;
        weights[ 687 ] <= 32'h bab07121 ;
        weights[ 688 ] <= 32'h b9b836cc ;
        weights[ 689 ] <= 32'h b7dc25dc ;
        weights[ 690 ] <= 32'h 384c2d85 ;
        weights[ 691 ] <= 32'h 389074b2 ;
        weights[ 692 ] <= 32'h 390406a4 ;
        weights[ 693 ] <= 32'h 38fb433a ;
        weights[ 694 ] <= 32'h 38bb9cb0 ;
        weights[ 695 ] <= 32'h 3761ce50 ;
        weights[ 696 ] <= 32'h b60d0ac5 ;
        weights[ 697 ] <= 32'h b628b925 ;
        weights[ 698 ] <= 32'h 353344b7 ;
        weights[ 699 ] <= 32'h 34bdd04a ;
        weights[ 700 ] <= 32'h 0 ;
        weights[ 701 ] <= 32'h 0 ;
        weights[ 702 ] <= 32'h 0 ;
        weights[ 703 ] <= 32'h 0 ;
        weights[ 704 ] <= 32'h 0 ;
        weights[ 705 ] <= 32'h 0 ;
        weights[ 706 ] <= 32'h 35d82d37 ;
        weights[ 707 ] <= 32'h 36827f33 ;
        weights[ 708 ] <= 32'h 36a8b927 ;
        weights[ 709 ] <= 32'h 374c5035 ;
        weights[ 710 ] <= 32'h 36a17932 ;
        weights[ 711 ] <= 32'h b800230d ;
        weights[ 712 ] <= 32'h b9910253 ;
        weights[ 713 ] <= 32'h 3a3e2f41 ;
        weights[ 714 ] <= 32'h 39b3a30a ;
        weights[ 715 ] <= 32'h 390dc2a1 ;
        weights[ 716 ] <= 32'h 38bd7cc6 ;
        weights[ 717 ] <= 32'h 378e5551 ;
        weights[ 718 ] <= 32'h 34d2e76e ;
        weights[ 719 ] <= 32'h b5812dc0 ;
        weights[ 720 ] <= 32'h 0 ;
        weights[ 721 ] <= 32'h 0 ;
        weights[ 722 ] <= 32'h 0 ;
        weights[ 723 ] <= 32'h 0 ;
        weights[ 724 ] <= 32'h 0 ;
        weights[ 725 ] <= 32'h 0 ;
        weights[ 726 ] <= 32'h 0 ;
        weights[ 727 ] <= 32'h 0 ;
        weights[ 728 ] <= 32'h 0 ;
        weights[ 729 ] <= 32'h 0 ;
        weights[ 730 ] <= 32'h 0 ;
        weights[ 731 ] <= 32'h 0 ;
        weights[ 732 ] <= 32'h 0 ;
        weights[ 733 ] <= 32'h 0 ;
        weights[ 734 ] <= 32'h 0 ;
        weights[ 735 ] <= 32'h 0 ;
        weights[ 736 ] <= 32'h 0 ;
        weights[ 737 ] <= 32'h 0 ;
        weights[ 738 ] <= 32'h 0 ;
        weights[ 739 ] <= 32'h 35c31613 ;
        weights[ 740 ] <= 32'h 355d7301 ;
        weights[ 741 ] <= 32'h 0 ;
        weights[ 742 ] <= 32'h 0 ;
        weights[ 743 ] <= 32'h 36e8f70c ;
        weights[ 744 ] <= 32'h 37add052 ;
        weights[ 745 ] <= 32'h 36e8f70c ;
        weights[ 746 ] <= 32'h 0 ;
        weights[ 747 ] <= 32'h 0 ;
        weights[ 748 ] <= 32'h 0 ;
        weights[ 749 ] <= 32'h 0 ;
        weights[ 750 ] <= 32'h 0 ;
        weights[ 751 ] <= 32'h 0 ;
        weights[ 752 ] <= 32'h 0 ;
        weights[ 753 ] <= 32'h 0 ;
        weights[ 754 ] <= 32'h 0 ;
        weights[ 755 ] <= 32'h 0 ;
        weights[ 756 ] <= 32'h 0 ;
        weights[ 757 ] <= 32'h 0 ;
        weights[ 758 ] <= 32'h 0 ;
        weights[ 759 ] <= 32'h 0 ;
        weights[ 760 ] <= 32'h 0 ;
        weights[ 761 ] <= 32'h 0 ;
        weights[ 762 ] <= 32'h 0 ;
        weights[ 763 ] <= 32'h 0 ;
        weights[ 764 ] <= 32'h 0 ;
        weights[ 765 ] <= 32'h 0 ;
        weights[ 766 ] <= 32'h 0 ;
        weights[ 767 ] <= 32'h 0 ;
        weights[ 768 ] <= 32'h 0 ;
        weights[ 769 ] <= 32'h 0 ;
        weights[ 770 ] <= 32'h 0 ;
        weights[ 771 ] <= 32'h 0 ;
        weights[ 772 ] <= 32'h 0 ;
        weights[ 773 ] <= 32'h 0 ;
        weights[ 774 ] <= 32'h 0 ;
        weights[ 775 ] <= 32'h 0 ;
        weights[ 776 ] <= 32'h 0 ;
        weights[ 777 ] <= 32'h 0 ;
        weights[ 778 ] <= 32'h 0 ;
        weights[ 779 ] <= 32'h 0 ;
        weights[ 780 ] <= 32'h 0 ;
        weights[ 781 ] <= 32'h 0 ;
        weights[ 782 ] <= 32'h 0 ;
        weights[ 783 ] <= 32'h 0 ;
        weights[ 784 ] <= 32'h 0 ;
		  data_out <= weights[addr];

		end
		else begin

			if (addr <= 10'd784)
				data_out <= weights[addr];
			else
				data_out <= 32'd0;
		end
	end
endmodule
